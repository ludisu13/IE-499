module wishbone (
	

);


endmodule
