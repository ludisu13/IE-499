module WB_(
input request,

ack,
writeread




);
