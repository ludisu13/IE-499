module cmd_controller(









);









endmodule 
